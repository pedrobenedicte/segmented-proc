LIBRARY ieee;
use ieee.std_logic_1164.all;
use IEEE.numeric_std.all;
use ieee.std_logic_unsigned.all;

entity ff_alu_lookup is 

end ff_alu_lookup;


architecture Structure of ff_alu_lookup is

begin


end Structure;