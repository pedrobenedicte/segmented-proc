LIBRARY ieee;
use ieee.std_logic_1164.all;
use IEEE.numeric_std.all;
use ieee.std_logic_unsigned.all;

entity stage_fwb is

end stage_fwb;


architecture Structure of stage_fwb is

begin


end Structure;
