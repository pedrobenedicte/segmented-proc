LIBRARY ieee;
use ieee.std_logic_1164.all;
use IEEE.numeric_std.all;
use ieee.std_logic_unsigned.all;

entity ff_fetch_decode is 

end ff_fetch_decode;


architecture Structure of ff_fetch_decode is

begin


end Structure;