// Module with global variables that will
// be used in the project

module global;

parameter NUM_BITS = 16;
parameter LOG_NUM_BITS = 4;

endmodule
