LIBRARY ieee;
use ieee.std_logic_1164.all;
use IEEE.numeric_std.all;
use ieee.std_logic_unsigned.all;

entity stage_wb is

end stage_wb;


architecture Structure of stage_wb is

begin


end Structure;
