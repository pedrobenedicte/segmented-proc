LIBRARY ieee;
USE ieee.std_logic_1164.all;
use IEEE.numeric_std.all;
USE ieee.std_logic_unsigned.all;

ENTITY ff_decode_alu IS 

END ff_decode_alu;


ARCHITECTURE Structure OF ff_decode_alu IS

BEGIN


END Structure;