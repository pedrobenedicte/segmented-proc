LIBRARY ieee;
use ieee.std_logic_1164.all;
use IEEE.numeric_std.all;
use ieee.std_logic_unsigned.all;

entity stage_fetch is

end stage_fetch;


architecture Structure of stage_fetch is

begin


end Structure;