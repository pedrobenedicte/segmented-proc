LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY proc IS

END proc;


ARCHITECTURE Structure OF proc IS

	COMPONENT datapath IS
	END COMPONENT;

	COMPONENT control_unit IS
	END COMPONENT;

BEGIN


END Structure;