LIBRARY ieee;
use ieee.std_logic_1164.all;
use IEEE.numeric_std.all;
use ieee.std_logic_unsigned.all;

entity stage_alu is

end stage_alu;


architecture Structure of stage_alu is

begin


end Structure;