LIBRARY ieee;
use ieee.std_logic_1164.all;
use IEEE.numeric_std.all;
use ieee.std_logic_unsigned.all;

entity stage_cache is

end stage_cache;


architecture Structure of stage_cache is

begin


end Structure;