LIBRARY ieee;
use ieee.std_logic_1164.all;
use IEEE.numeric_std.all;
use ieee.std_logic_unsigned.all;

entity ff_lookup_cache is 

end ff_lookup_cache;


architecture Structure of ff_lookup_cache is

begin


end Structure;