LIBRARY ieee;
use ieee.std_logic_1164.all;
use IEEE.numeric_std.all;
use ieee.std_logic_unsigned.all;

entity stage_lookup is

end stage_lookup;


architecture Structure of stage_lookup is

begin


end Structure;