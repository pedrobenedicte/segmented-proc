LIBRARY ieee;
USE ieee.std_logic_1164.all;

entity proc is

end proc;


architecture Structure of proc is

	component datapath is
	end component;

	component control_unit is
	end component;

begin


end Structure;