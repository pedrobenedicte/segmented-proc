LIBRARY ieee;
USE ieee.std_logic_1164.all;
use IEEE.numeric_std.all;
USE ieee.std_logic_unsigned.all;

ENTITY control_unit IS 

END control_unit;


ARCHITECTURE Structure OF control_unit IS

BEGIN


END Structure;