LIBRARY ieee;
use ieee.std_logic_1164.all;
use IEEE.numeric_std.all;
use ieee.std_logic_unsigned.all;

entity ff_f5_fwb is 

end ff_f5_fwb;


architecture Structure of ff_f5_fwb is

begin


end Structure;
