LIBRARY ieee;
use ieee.std_logic_1164.all;
use IEEE.numeric_std.all;
use ieee.std_logic_unsigned.all;

entity ff_cache_wb is 
	port (
		clk			: in	std_logic;
		stall		: in	std_logic;
		nop			: in	std_logic
	);
end ff_cache_wb;


architecture Structure of ff_cache_wb is

begin


end Structure;