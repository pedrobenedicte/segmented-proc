LIBRARY ieee;
use ieee.std_logic_1164.all;
use IEEE.numeric_std.all;
use ieee.std_logic_unsigned.all;

entity stage_decode is

end stage_decode;


architecture Structure of stage_decode is

begin


end Structure;