LIBRARY ieee;
use ieee.std_logic_1164.all;
use IEEE.numeric_std.all;
use ieee.std_logic_unsigned.all;

entity stage_f5 is

end stage_f5;


architecture Structure of stage_f5 is

begin


end Structure;
