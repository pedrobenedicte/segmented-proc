LIBRARY ieee;
use ieee.std_logic_1164.all;
use IEEE.numeric_std.all;
use ieee.std_logic_unsigned.all;

entity ff_decode_alu is 

end ff_decode_alu;


architecture Structure of ff_decode_alu is

begin


end Structure;