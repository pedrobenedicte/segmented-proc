// 

module adder(input [15:0] A, input [15:0] B, output cout, output [15:0] sum);

wire 

endmodule
