LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY test_proc IS 


END test_proc;


ARCHITECTURE Structure OF test_proc IS


BEGIN


END Structure;