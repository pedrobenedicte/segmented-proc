LIBRARY ieee;
use ieee.std_logic_1164.all;
use IEEE.numeric_std.all;
use ieee.std_logic_unsigned.all;

entity stage_fwb is
	port (
		clk			: in	std_logic;
		rdest		: in	std_logic_vector(2 downto 0)
	);
end stage_fwb;


architecture Structure of stage_fwb is

begin


end Structure;
