LIBRARY ieee;
USE ieee.std_logic_1164.all;
use IEEE.numeric_std.all;
USE ieee.std_logic_unsigned.all;

ENTITY datapath IS 

END datapath;


ARCHITECTURE Structure OF datapath IS

BEGIN

	-- Stages and interconnection between stages

END Structure;