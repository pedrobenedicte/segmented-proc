LIBRARY ieee;
USE ieee.std_logic_1164.all;
use IEEE.numeric_std.all;
USE ieee.std_logic_unsigned.all;

ENTITY stage_decode IS 

END stage_decode;


ARCHITECTURE Structure OF stage_decode IS

BEGIN


END Structure;